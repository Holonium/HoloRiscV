/*

This version of the core is designed for implementation on a chip. Currently, only the RV32I ISA is being implemented.
The exception to this is the EBREAK, ECALL, and FENCE instructions.
The pipeline is composed of 5 stages, none of which currently run in parallel.

*/

`default_nettype none

module HoloRiscV (

	);
	
endmodule
